module led2sw(output led_o, input sw_i);

assign led_o = sw_i;

endmodule