module ex3();

endmodule