`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:13:59 03/04/2019 
// Design Name: 
// Module Name:    MY_XOR_3 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module MY_XOR_3(
    input A,
    input B,
    input C,
    output O
    );

assign 0 = A^B^C;
endmodule
