`timescale 1 ns/1 ps
module hex_7display
(input [3:0] c,
output [6:0] hex,
output cut
);
assign cut = 1;
assign hex[0] = ~((~c[2]&~c[0])|(~c[3]&c[1])|(~c[3]&c[2]&c[0])|(c[3]&~c[2]&~c[1])|(c[3]&~c[0])|(c[2]&c[1]));//A
assign hex[1] = ~((~c[2]&~c[0])|(~c[3]&~c[2])|(c[3]&~c[1]&c[0])|(~c[3]&c[1]&c[0])|(~c[3]&~c[1]&~c[0])); //B
assign hex[2] = ~((c[3]&~c[2])|(~c[3]&c[2])|(~c[1]&c[0])|(~c[3]&~c[2]&~c[1])|(~c[3]&~c[2]&c[0])); //C
assign hex[3] = ~((c[3]&~c[1]&~c[0])|(c[2]&~c[1]&c[0])|(~c[2]&c[1]&c[0])|(c[2]&c[1]&~c[0])|(~c[3]&~c[2]&~c[0]));//D
assign hex[4] = ~((~c[2]&~c[0])|(c[3]&c[2])|(c[1]&~c[0])|(c[3]&c[1]));//E
assign hex[5] = ~((~c[1]&~c[0])|(c[3]&~c[2])|(c[3]&c[1])|(~c[3]&c[2]&~c[1])|(~c[3]&c[2]&~c[0])); //F
assign hex[6] = ~((c[1]&~c[0])|(c[3]&~c[2])|(c[3]&c[0])|(~c[3]&c[2]&~c[1])|(~c[3]&~c[2]&c[1]));//G
 endmodule