module main;

initial 
	$display("Hello, world!");
//pentru run do run_helloWorld.txt
//vsim -topargs ---> pune numele modulului
//iar la catch numele fisierului
endmodule
